

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO System_Top 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 0.241 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.15921 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 27.774 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 133.785 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 628.605 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3037.38 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 0.291 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.39971 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.14862 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 26.708 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 128.658 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 577.025 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2785.37 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 4.843 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2948 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.97 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4805 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 82.8077 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 408.483 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.3546 LAYER VIA34 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 2.089 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2405 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 41.8133 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 204.081 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.677298 LAYER VIA23 ;
  END SI[0]
  PIN SO[3] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.854 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.1625 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 59.5819 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 285.135 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.20736 LAYER VIA34 ;
  END SO[3]
  PIN SO[2] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.177 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.85377 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 35.048 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 168.966 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4563 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 128.291 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 624.061 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.93337 LAYER VIA56 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.679 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.45839 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 29.824 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 143.646 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 158.201 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 764.35 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.09372 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 1.815 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.92255 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 16.685 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 80.6397 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 277.915 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1346.81 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.4868 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 22.362 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 107.754 LAYER METAL5 ;
    ANTENNAGATEAREA 0.3133 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 349.291 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1690.74 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.4868 LAYER VIA56 ;
  END SO[0]
  PIN SE 
    ANTENNAPARTIALMETALAREA 0.273 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.31313 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 7.77379 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 35.0467 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.205698 LAYER VIA23 ;
  END SE
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.255 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.22655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.124 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59884 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.99326 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 1.53833 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 7.54512 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 0.223 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.07263 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.42 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6426 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 7.337 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.6758 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 7.086 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.4685 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 85.7599 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 418.665 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.551 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.65031 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 17.9036 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 89.5299 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.828932 LAYER VIA34 ;
  END test_mode
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.291 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.39971 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 3.8408 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 18.62 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END REF_CLK
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.487 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.34247 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.994 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.4035 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 1.46422 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 7.12581 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END UART_CLK
  PIN RST 
    ANTENNAPARTIALMETALAREA 0.893 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.29533 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.14862 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 69.8124 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 339.551 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.3546 LAYER VIA34 ;
  END RST
  PIN RX_IN 
    ANTENNAPARTIALMETALAREA 0.997 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.79557 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04906 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 14.326 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 69.1005 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6552 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 48.3565 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 235.057 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.4243 LAYER VIA56 ;
  END RX_IN
  PIN Stop_Error 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.194 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL3 ;
  END Stop_Error
  PIN Parity_Error 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.527 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1573 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 26.38 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 127.08 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3406 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 110.345 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 533.407 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.56658 LAYER VIA56 ;
  END Parity_Error
  PIN TX_OUT 
    ANTENNADIFFAREA 0.952 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.998 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.61038 LAYER METAL3 ;
  END TX_OUT
END System_Top

END LIBRARY
